library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package custom_flow is
	   type COLOR_DATA is array(0 to 2) of std_logic_vector(9 downto 0);
	   type COLOR is array(0 to 11) of COLOR_DATA; 
	   constant data : COLOR := (
 	   --(R,G,B)
	   ("0000000000","1111111100","1111111100"), --aqua blue
	   ("0000000000","0000000000","1111111100"), --regular blue
	   ("1000101100","0000000000","0000000000"), --dark red
	   ("0000000000","1000000000","0000000000"), --green
	   ("1111111100","1111111100","0000000000"), --yellow
	   ("1111111100","0000000000","0000000000"), --red
	   ("1000000000","0000000000","1000000000"), --purple
	   ("1111111100","1100000000","1100101100"), --pink
	   ("1111111100","1010010100","0000000000"), --orange
	   ("0000000000","1111111100","0000000000"), --lime
	   ("0000000000","1000000000","1000000000"), --teal
	   ("1000000000","1000000000","1000000000")  --gray
 	   ); 

 	   	type REG is array (0 to 35) of std_logic_vector(9 downto 0);
 	   	
 	   	--convention used here: 0 -> x_coord, 1 -> y_coord
	   type BLOCKS is array (0 to 11) of std_logic_vector(9 downto 0);
	   type COLOR_TYPE is array (0 to 11) of integer range 0 to 11;
	   type COORDS is array (0 to 11) of integer range 0 to 35;
	   type DATA_UNIT is array (0 to 144) of std_logic_vector(9 downto 0);


	   constant BOX_WIDTH: integer := 40;
	   constant BOX_HEIGHT: integer := 40;
	   constant Step    : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(40, 10);  --Leftmost point on the X axis
	   constant X_Min    : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(80, 10);  --Leftmost point on the X axis
	   constant X_Max    : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(560, 10);  --Rightmost point on the X axis
	   constant Y_Min    : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(0, 10);   --Topmost point on the Y axis
	   constant Y_Max    : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(480, 10);  --Bottommost point on the Y axis
	   
	   
	   -- level 21 on iphone game
	   constant blk0_x : BLOCKS := ("0100011000","0001111000","0100011000","0110010000","0001111000","0010100000",
									"0110111000","0101000000","0011110000","0011001000","0101000000","1010000000"); 
	   constant blk1_x : BLOCKS := ("0110010000","0101000000","0110010000","0111100000","0010100000","0001111000",
									"0110111000","0011110000","0111100000","0010100000","0110010000","1010000000");
		constant blk0_y : BLOCKS := ("0000000000","0000101000","0000101000","0000101000","0001010000","0001010000",
									"0001010000","0010100000","0011110000","0100011000","0101101000","1010000000");
	   constant blk1_y : BLOCKS := ("0110010000","0001010000","0011001000","0101101000","0011001000","0110010000",
									"0011001000","0101101000","0110010000","0110010000","0101101000","1010000000");
		-- level 22 on iphone game
									
									
--		constant blk0_x : BLOCKS := ("0001111000", "0010100000", "0110010000", "0001010000", "0101000000", "0001111000",
--									"0010100000", "0101000000", "0010100000", "0110010000", "0101000000", "1010000000");
--		constant blk0_y : BLOCKS := ( "0000101000", "0000101000", "0001111000", "0010100000", "0010100000", "0011110000",
--									"0011110000", "0011110000", "0100011000", "0100011000", "0101000000", "1010000000");				
--		constant blk1_y : BLOCKS := ("0011110000", "0100011000", "0101101000", "0010100000", "0100011000", "0010100000",
--									"0011110000", "0010100000", "0001010000", "0100011000", "0110010000", "1010000000");
--		constant blk1_x : BLOCKS := ("0011110000","0100011000","0101101000","0010100000","0100011000","0010100000",
--									"0011110000","0010100000","0001010000","0100011000","0110010000","1010000000");	
										
				
   constant ADDR_WIDTH: integer:=11;
   constant DATA_WIDTH: integer:=8;
   type rom_type is array (0 to 95)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant ROM: rom_type:=(
   
   "00000000", -- 0
   "00000000", -- 1
   "11000011", -- 2 **    **
   "11000011", -- 3 **    **
   "11000011", -- 4 **    **
   "01100110", -- 5  **  **
   "00111100", -- 6   ****
   "00011000", -- 7    **
   "00011000", -- 8    **
   "00011000", -- 9    **
   "00011000", -- a    **
   "00111100", -- b   ****
   "00000000", -- c
   "00000000", -- d
   "00000000", -- e
   "00000000", -- f

   "00000000", -- 0
   "00000000", -- 1
   "01111100", -- 2  *****
   "11000110", -- 3 **   **
   "11000110", -- 4 **   **
   "11000110", -- 5 **   **
   "11000110", -- 6 **   **
   "11000110", -- 7 **   **
   "11000110", -- 8 **   **
   "11000110", -- 9 **   **
   "11000110", -- a **   **
   "01111100", -- b  *****
   "00000000", -- c
   "00000000", -- d
   "00000000", -- e
   "00000000", -- f

   "00000000", -- 0
   "00000000", -- 1
   "11000110", -- 2 **   **
   "11000110", -- 3 **   **
   "11000110", -- 4 **   **
   "11000110", -- 5 **   **
   "11000110", -- 6 **   **
   "11000110", -- 7 **   **
   "11000110", -- 8 **   **
   "11000110", -- 9 **   **
   "11000110", -- a **   **
   "01111100", -- b  *****
   "00000000", -- c
   "00000000", -- d
   "00000000", -- e
   "00000000", -- f

   "00000000", -- 0
   "00000000", -- 1
   "11000011", -- 2 **    **
   "11000011", -- 3 **    **
   "11000011", -- 4 **    **
   "11000011", -- 5 **    **
   "11000011", -- 6 **    **
   "11011011", -- 7 ** ** **
   "11011011", -- 8 ** ** **
   "11111111", -- 9 ********
   "01100110", -- a  **  **
   "01100110", -- b  **  **
   "00000000", -- c
   "00000000", -- d
   "00000000", -- e
   "00000000", -- f

   "00000000", -- 0
   "00000000", -- 1
   "00111100", -- 2   ****
   "00011000", -- 3    **
   "00011000", -- 4    **
   "00011000", -- 5    **
   "00011000", -- 6    **
   "00011000", -- 7    **
   "00011000", -- 8    **
   "00011000", -- 9    **
   "00011000", -- a    **
   "00111100", -- b   ****
   "00000000", -- c
   "00000000", -- d
   "00000000", -- e
   "00000000", -- f


   "00000000", -- 0
   "00000000", -- 1
   "11000110", -- 2 **   **
   "11100110", -- 3 ***  **
   "11110110", -- 4 **** **
   "11111110", -- 5 *******
   "11011110", -- 6 ** ****
   "11001110", -- 7 **  ***
   "11000110", -- 8 **   **
   "11000110", -- 9 **   **
   "11000110", -- a **   **
   "11000110", -- b **   **
   "00000000", -- c
   "00000000", -- d
   "00000000", -- e
   "00000000" -- f
   
   );
	   
   
end custom_flow;

package body custom_flow is
     -- Definition of previously declared
        -- constants
        -- subprograms
     -- Declaration/definition of additional
        -- types and subtypes
        -- subprograms
        -- constants, signals and shared variables
end custom_flow;